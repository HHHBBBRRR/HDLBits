module top_module (
	input clk,
	input L,
	input r_in,
	input q_in,
	output reg Q
);
    wire wire1;

    assign wire1 = L ? r_in : q_in;

    always @(posedge clk) begin
        Q <= wire1;
    end

endmodule
